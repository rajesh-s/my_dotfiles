//https://www.veripool.org/projects/verilog-mode/wiki/Faq
module samp;
pinmux_top pmux (
/*AUTOINST*/
endmodule
// Local Variables:
// verilog-library-directories:(".")
// End:
